
entity normalization_controller is
end normalization_controller;
