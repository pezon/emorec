library ieee;

entity chisquare_tb is
end chisquare_tb;

architecture tb of chisquare_tb is
begin
end tb;

