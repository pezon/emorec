library ieee;

use ieee.std_logic_1164.all;

entity emorec_datapath is
end emorec_datapath;

