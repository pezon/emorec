library ieee;

use ieee.std_logic_1164.all;

entity emorec_controller is
end emorec_controller;

