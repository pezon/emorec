
entity chisquare_controller is
end chisquare_controller;
