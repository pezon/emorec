library ieee;

use ieee.std_logic_1164.all;

entity top_level is
end top_level;

